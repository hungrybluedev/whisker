module whisker
